`timescale 1nd/1ns

module IF_Stage 
(
    input clk, rst, branch_taken,
    input [31:0] BranchAddr,
    output [31:0] PC, Instruction
);



    
endmodule