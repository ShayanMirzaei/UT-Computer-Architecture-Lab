`timescale 1nd/1ns

module IF_Stage_Register
(
    input clk, rst, freeze, flush
    input [31:0] PC_in, Instruction_in,
    output reg [31:0] PC, Instruction
);



    
endmodule