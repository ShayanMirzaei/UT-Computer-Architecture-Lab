`timescale 1nd/1ns

module EXE_Stage_Reg
(
    input clk, rst,
    input [31:0] PC_in,
    output reg [31:0] PC
);



    
endmodule